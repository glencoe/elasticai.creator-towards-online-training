entity ${name} is
end;

architecture rtl of ${name} is

begin
end;